module multiplicador_uc(
     input  clk, rst, start, qlsb, zero,
     output a_rst, a_en, b_en, q_en, cnt_en,
            a_ld, b_ld, q_ld, cnt_ld, done
);


endmodule